module example(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h0c000003;
30'h00000002: inst = 32'h37bd0100;
30'h00000003: inst = 32'h27bdffe0;
30'h00000004: inst = 32'hafbe0018;
30'h00000005: inst = 32'h03a0f021;
30'h00000006: inst = 32'h24020064;
30'h00000007: inst = 32'hafc20014;
30'h00000008: inst = 32'h8fc20014;
30'h00000009: inst = 32'h00000000;
30'h0000000a: inst = 32'h244201f4;
30'h0000000b: inst = 32'hafc20010;
30'h0000000c: inst = 32'h240203e8;
30'h0000000d: inst = 32'hafc2000c;
30'h0000000e: inst = 32'h8fc2000c;
30'h0000000f: inst = 32'h00000000;
30'h00000010: inst = 32'h00021027;
30'h00000011: inst = 32'hafc20008;
30'h00000012: inst = 32'h3c021000;
30'h00000013: inst = 32'h2442011c;
30'h00000014: inst = 32'h90420003;
30'h00000015: inst = 32'h00000000;
30'h00000016: inst = 32'ha3c20004;
30'h00000017: inst = 32'h3c021000;
30'h00000018: inst = 32'h2443011c;
30'h00000019: inst = 32'h24020042;
30'h0000001a: inst = 32'ha0620004;
30'h0000001b: inst = 32'h3c021000;
30'h0000001c: inst = 32'h2443011c;
30'h0000001d: inst = 32'h24020043;
30'h0000001e: inst = 32'ha0620005;
30'h0000001f: inst = 32'h3c021000;
30'h00000020: inst = 32'h2443011c;
30'h00000021: inst = 32'h24020044;
30'h00000022: inst = 32'ha0620006;
30'h00000023: inst = 32'h3c021000;
30'h00000024: inst = 32'h2443011c;
30'h00000025: inst = 32'h24020045;
30'h00000026: inst = 32'ha0620007;
30'h00000027: inst = 32'h3c021000;
30'h00000028: inst = 32'h2442011c;
30'h00000029: inst = 32'h90420004;
30'h0000002a: inst = 32'h00000000;
30'h0000002b: inst = 32'ha3c20003;
30'h0000002c: inst = 32'h3c021000;
30'h0000002d: inst = 32'h2442011c;
30'h0000002e: inst = 32'h90420005;
30'h0000002f: inst = 32'h00000000;
30'h00000030: inst = 32'ha3c20002;
30'h00000031: inst = 32'h3c021000;
30'h00000032: inst = 32'h2442011c;
30'h00000033: inst = 32'h90420006;
30'h00000034: inst = 32'h00000000;
30'h00000035: inst = 32'ha3c20001;
30'h00000036: inst = 32'h3c021000;
30'h00000037: inst = 32'h2442011c;
30'h00000038: inst = 32'h90420007;
30'h00000039: inst = 32'h00000000;
30'h0000003a: inst = 32'ha3c20000;
30'h0000003b: inst = 32'h8fc20010;
30'h0000003c: inst = 32'h03c0e821;
30'h0000003d: inst = 32'h8fbe0018;
30'h0000003e: inst = 32'h27bd0020;
30'h0000003f: inst = 32'h03e00008;
30'h00000040: inst = 32'h00000000;
30'h00000041: inst = 32'h00000003;
30'h00000042: inst = 32'h00000002;
30'h00000043: inst = 32'h00000004;
30'h00000044: inst = 32'h00000017;
30'h00000045: inst = 32'h00000020;
30'h00000046: inst = 32'h00000001;
30'h00000047: inst = 32'h48454c4c;
30'h00000048: inst = 32'h4f20574f;
30'h00000049: inst = 32'h524c4421;
30'h0000004a: inst = 32'h21000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
